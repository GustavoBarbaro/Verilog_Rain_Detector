module Memoria_Mensagem (input [2:0] flag_mensagem,

		output reg [7:0] hex_1_00, hex_1_01, hex_1_02, hex_1_03, hex_1_04, hex_1_05, hex_1_06, hex_1_07, hex_1_08, hex_1_09, hex_1_10, hex_1_11, hex_1_12, hex_1_13, hex_1_14, hex_1_15,
		output reg [7:0] hex_2_00, hex_2_01, hex_2_02, hex_2_03, hex_2_04, hex_2_05, hex_2_06, hex_2_07, hex_2_08, hex_2_09, hex_2_10, hex_2_11, hex_2_12, hex_2_13, hex_2_14, hex_2_15


);






	always @ (flag_mensagem) begin
	
	
	// se enable = 1 entao pode escrever chovendo/ seco etc
	//se for 0 então é display limpo

		case (flag_mensagem)
		
			3'b000: begin //display limpo
			
				hex_1_00 = 8'h00000020;
				hex_1_01 = 8'h00000020;
				hex_1_02 = 8'h00000020;
				hex_1_03 = 8'h00000020;
				hex_1_04 = 8'h00000020;
				hex_1_05 = 8'h00000020;
				hex_1_06 = 8'h00000020;
				hex_1_07 = 8'h00000020;
				hex_1_08 = 8'h00000020;
				hex_1_09 = 8'h00000020;
				hex_1_10 = 8'h00000020;
				hex_1_11 = 8'h00000020;
				hex_1_12 = 8'h00000020;
				hex_1_13 = 8'h00000020;
				hex_1_14 = 8'h00000020;
				hex_1_15 = 8'h00000020;
				
				hex_2_00 = 8'h00000020;
				hex_2_01 = 8'h00000020;
				hex_2_02 = 8'h00000020;
				hex_2_03 = 8'h00000020;
				hex_2_04 = 8'h00000020;
				hex_2_05 = 8'h00000020;
				hex_2_06 = 8'h00000020;
				hex_2_07 = 8'h00000020;
				hex_2_08 = 8'h00000020;
				hex_2_09 = 8'h00000020;
				hex_2_10 = 8'h00000020;
				hex_2_11 = 8'h00000020;
				hex_2_12 = 8'h00000020;
				hex_2_13 = 8'h00000020;
				hex_2_14 = 8'h00000020;
				hex_2_15 = 8'h00000020;
			
			end
		
		
			3'b001: begin //Chovendo !
			
				hex_1_00 = 8'h00000043;
				hex_1_01 = 8'h00000068;
				hex_1_02 = 8'h0000006f;
				hex_1_03 = 8'h00000076;
				hex_1_04 = 8'h00000065;
				hex_1_05 = 8'h0000006e;
				hex_1_06 = 8'h00000064;
				hex_1_07 = 8'h0000006f;
				hex_1_08 = 8'h00000020;
				hex_1_09 = 8'h00000021;
				hex_1_10 = 8'h00000020;
				hex_1_11 = 8'h00000020;
				hex_1_12 = 8'h00000020;
				hex_1_13 = 8'h00000020;
				hex_1_14 = 8'h00000020;
				hex_1_15 = 8'h00000020;

				hex_2_00 = 8'h00000020;
				hex_2_01 = 8'h00000020;
				hex_2_02 = 8'h00000020;
				hex_2_03 = 8'h00000020;
				hex_2_04 = 8'h00000020;
				hex_2_05 = 8'h00000020;
				hex_2_06 = 8'h00000020;
				hex_2_07 = 8'h00000020;
				hex_2_08 = 8'h00000020;
				hex_2_09 = 8'h00000020;
				hex_2_10 = 8'h00000020;
				hex_2_11 = 8'h00000020;
				hex_2_12 = 8'h00000020;
				hex_2_13 = 8'h00000020;
				hex_2_14 = 8'h00000020;
				hex_2_15 = 8'h00000020;
			
			end
			
			
			3'b010: begin // Tempo seco !
			
				hex_1_00 = 8'h00000054;
				hex_1_01 = 8'h00000065;
				hex_1_02 = 8'h0000006d;
				hex_1_03 = 8'h00000070;
				hex_1_04 = 8'h0000006f;
				hex_1_05 = 8'h00000020;
				hex_1_06 = 8'h00000053;
				hex_1_07 = 8'h00000065;
				hex_1_08 = 8'h00000063;
				hex_1_09 = 8'h0000006f;
				hex_1_10 = 8'h00000020;
				hex_1_11 = 8'h00000021;
				hex_1_12 = 8'h00000020;
				hex_1_13 = 8'h00000020;
				hex_1_14 = 8'h00000020;
				hex_1_15 = 8'h00000020;

				hex_2_00 = 8'h00000020;
				hex_2_01 = 8'h00000020;
				hex_2_02 = 8'h00000020;
				hex_2_03 = 8'h00000020;
				hex_2_04 = 8'h00000020;
				hex_2_05 = 8'h00000020;
				hex_2_06 = 8'h00000020;
				hex_2_07 = 8'h00000020;
				hex_2_08 = 8'h00000020;
				hex_2_09 = 8'h00000020;
				hex_2_10 = 8'h00000020;
				hex_2_11 = 8'h00000020;
				hex_2_12 = 8'h00000020;
				hex_2_13 = 8'h00000020;
				hex_2_14 = 8'h00000020;
				hex_2_15 = 8'h00000020;
			
			end
			
			3'b011: begin // Bluetooth on
			
				hex_1_00 = 8'h00000042;
				hex_1_01 = 8'h0000006c;
				hex_1_02 = 8'h00000075;
				hex_1_03 = 8'h00000065;
				hex_1_04 = 8'h00000074;
				hex_1_05 = 8'h0000006f;
				hex_1_06 = 8'h0000006f;
				hex_1_07 = 8'h00000074;
				hex_1_08 = 8'h00000068;
				hex_1_09 = 8'h0000003a;
				hex_1_10 = 8'h00000020;
				hex_1_11 = 8'h00000020;
				hex_1_12 = 8'h00000020;
				hex_1_13 = 8'h00000020;
				hex_1_14 = 8'h00000020;
				hex_1_15 = 8'h00000020;

				hex_2_00 = 8'h0000004f;
				hex_2_01 = 8'h0000006e;
				hex_2_02 = 8'h00000020;
				hex_2_03 = 8'h00000020;
				hex_2_04 = 8'h00000020;
				hex_2_05 = 8'h00000020;
				hex_2_06 = 8'h00000020;
				hex_2_07 = 8'h00000020;
				hex_2_08 = 8'h00000020;
				hex_2_09 = 8'h00000020;
				hex_2_10 = 8'h00000020;
				hex_2_11 = 8'h00000020;
				hex_2_12 = 8'h00000020;
				hex_2_13 = 8'h00000020;
				hex_2_14 = 8'h00000020;
				hex_2_15 = 8'h00000020;
			
			end
			
			
			3'b100: begin // Bluetooth off
			
				hex_1_00 = 8'h00000042;
				hex_1_01 = 8'h0000006c;
				hex_1_02 = 8'h00000075;
				hex_1_03 = 8'h00000065;
				hex_1_04 = 8'h00000074;
				hex_1_05 = 8'h0000006f;
				hex_1_06 = 8'h0000006f;
				hex_1_07 = 8'h00000074;
				hex_1_08 = 8'h00000068;
				hex_1_09 = 8'h0000003a;
				hex_1_10 = 8'h00000020;
				hex_1_11 = 8'h00000020;
				hex_1_12 = 8'h00000020;
				hex_1_13 = 8'h00000020;
				hex_1_14 = 8'h00000020;
				hex_1_15 = 8'h00000020;

				hex_2_00 = 8'h0000004f;
				hex_2_01 = 8'h00000066;
				hex_2_02 = 8'h00000066;
				hex_2_03 = 8'h00000020;
				hex_2_04 = 8'h00000020;
				hex_2_05 = 8'h00000020;
				hex_2_06 = 8'h00000020;
				hex_2_07 = 8'h00000020;
				hex_2_08 = 8'h00000020;
				hex_2_09 = 8'h00000020;
				hex_2_10 = 8'h00000020;
				hex_2_11 = 8'h00000020;
				hex_2_12 = 8'h00000020;
				hex_2_13 = 8'h00000020;
				hex_2_14 = 8'h00000020;
				hex_2_15 = 8'h00000020;
			
			end
			
			3'b101: begin // Sensor desligado //Bluetooth: Off
			
				hex_1_00 = 8'h00000053;
				hex_1_01 = 8'h00000065;
				hex_1_02 = 8'h0000006e;
				hex_1_03 = 8'h00000073;
				hex_1_04 = 8'h0000006f;
				hex_1_05 = 8'h00000072;
				hex_1_06 = 8'h00000020;
				hex_1_07 = 8'h00000064;
				hex_1_08 = 8'h00000065;
				hex_1_09 = 8'h00000073;
				hex_1_10 = 8'h0000006c;
				hex_1_11 = 8'h00000069;
				hex_1_12 = 8'h00000067;
				hex_1_13 = 8'h00000061;
				hex_1_14 = 8'h00000064;
				hex_1_15 = 8'h0000006f;

				hex_2_00 = 8'h00000042;
				hex_2_01 = 8'h0000006c;
				hex_2_02 = 8'h00000075;
				hex_2_03 = 8'h00000065;
				hex_2_04 = 8'h00000074;
				hex_2_05 = 8'h0000006f;
				hex_2_06 = 8'h0000006f;
				hex_2_07 = 8'h00000074;
				hex_2_08 = 8'h00000068;
				hex_2_09 = 8'h0000003a;
				hex_2_10 = 8'h00000020;
				hex_2_11 = 8'h0000004f;
				hex_2_12 = 8'h00000066;
				hex_2_13 = 8'h00000066;
				hex_2_14 = 8'h00000020;
				hex_2_15 = 8'h00000020;
			
			end
			
			3'b110: begin // Bluetooth Reset
			
				hex_1_00 = 8'h00000042;
				hex_1_01 = 8'h0000006c;
				hex_1_02 = 8'h00000075;
				hex_1_03 = 8'h00000065;
				hex_1_04 = 8'h00000074;
				hex_1_05 = 8'h0000006f;
				hex_1_06 = 8'h0000006f;
				hex_1_07 = 8'h00000074;
				hex_1_08 = 8'h00000068;
				hex_1_09 = 8'h0000003a;
				hex_1_10 = 8'h00000020;
				hex_1_11 = 8'h00000020;
				hex_1_12 = 8'h00000020;
				hex_1_13 = 8'h00000020;
				hex_1_14 = 8'h00000020;
				hex_1_15 = 8'h00000020;

				hex_2_00 = 8'h00000052;
				hex_2_01 = 8'h00000065;
				hex_2_02 = 8'h00000073;
				hex_2_03 = 8'h00000065;
				hex_2_04 = 8'h00000074;
				hex_2_05 = 8'h00000021;
				hex_2_06 = 8'h00000020;
				hex_2_07 = 8'h00000020;
				hex_2_08 = 8'h00000020;
				hex_2_09 = 8'h00000020;
				hex_2_10 = 8'h00000020;
				hex_2_11 = 8'h00000020;
				hex_2_12 = 8'h00000020;
				hex_2_13 = 8'h00000020;
				hex_2_14 = 8'h00000020;
				hex_2_15 = 8'h00000020;
			
			end
			
			default: begin //display limpo
				hex_1_00 = 8'h00000020;
				hex_1_01 = 8'h00000020;
				hex_1_02 = 8'h00000020;
				hex_1_03 = 8'h00000020;
				hex_1_04 = 8'h00000020;
				hex_1_05 = 8'h00000020;
				hex_1_06 = 8'h00000020;
				hex_1_07 = 8'h00000020;
				hex_1_08 = 8'h00000020;
				hex_1_09 = 8'h00000020;
				hex_1_10 = 8'h00000020;
				hex_1_11 = 8'h00000020;
				hex_1_12 = 8'h00000020;
				hex_1_13 = 8'h00000020;
				hex_1_14 = 8'h00000020;
				hex_1_15 = 8'h00000020;

				hex_2_00 = 8'h00000020;
				hex_2_01 = 8'h00000020;
				hex_2_02 = 8'h00000020;
				hex_2_03 = 8'h00000020;
				hex_2_04 = 8'h00000020;
				hex_2_05 = 8'h00000020;
				hex_2_06 = 8'h00000020;
				hex_2_07 = 8'h00000020;
				hex_2_08 = 8'h00000020;
				hex_2_09 = 8'h00000020;
				hex_2_10 = 8'h00000020;
				hex_2_11 = 8'h00000020;
				hex_2_12 = 8'h00000020;
				hex_2_13 = 8'h00000020;
				hex_2_14 = 8'h00000020;
				hex_2_15 = 8'h00000020;
			end
		
		
		endcase
	end



endmodule